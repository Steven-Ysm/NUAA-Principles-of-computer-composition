`include "./datapath/pc.v"
`include "./datapath/npc.v"
`include "./datapath/pc_add4.v"
`include "./datapath/im.v"
`include "./datapath/IF_ID.v"
`include "./datapath/registerfile.v"
`include "./datapath/ID_EX.v"
`include "./datapath/alu.v"
`include "./datapath/aluctrl.v"
`include "./datapath/EX_MEM.v"
`include "./datapath/dm.v"
`include "./datapath/MEM_WB.v"
`include "./datapath/ext.v"
`include "./datapath/mux.v"

module data_path (RegDst, Jump, Branch, MemRead, MemtoReg, ALUOp, 
    MemWrite, ALUSrc, RegWrite, ExtOp, clk, rst, ID_ins);
    
    input                  RegDst;
    input                  Jump;
    input                  Branch;
    input                  MemRead;
    input                  MemtoReg;
    input [2: 0] ALUOp;
    input                  MemWrite;
    input                  ALUSrc;
    input                  RegWrite;
    input                  ExtOp;

    input                  clk;
    input                  rst;

    output [31: 0]         ID_ins;

    //IF_ID
    wire    [31:0] ID_PC;
    wire    [31:0] ID_ins;

    //ID_EX
    wire           EX_MemtoReg;
    wire           EX_RegWrite;
    wire           EX_Branch;
    wire           EX_Jump;
    wire           EX_MemWrite;
    wire           EX_MemRead;
    wire           EX_RegDst;
    wire           EX_ALUSrc;
    wire           EX_ExtOp;
    wire    [2:0] EX_ALUOp;
    wire    [31:0] EX_PC;
    wire    [25:0] EX_Jump_ins_add;
    wire    [31:0] EX_Reg_data_1_out;
    wire    [31:0] EX_Reg_data_2_out;
    wire    [15:0] EX_Extimm;
    wire    [4:0]  EX_rt;
    wire    [4:0]  EX_rd;
    //EX_MEM
    wire           MEM_MemtoReg;
    wire           MEM_RegWrite;
    wire           MEM_Branch;
    wire           MEM_Jump;
    wire           MEM_MemWrite;
    wire           MEM_MemRead;
    wire    [31:0] MEM_PC;
    wire    [25:0] MEM_Jump_ins_add;
    wire           MEM_Zero;
    wire    [31:0] MEM_ALU;
    wire    [31:0] MEM_WriteData;
    wire    [31:0] MEM_Extimm;
    wire    [4:0]  MEM_Reg_Write;
    //MEM_WB
    wire           WB_MemtoReg;
    wire           WB_RegWrite;
    wire    [31:0] WB_Data_out;
    wire    [31:0] WB_ALU;
    wire    [4:0]  WB_Reg_Write;

    // module wire
    wire    [31: 0] PC;             // value of pc
    wire    [31: 0] PC_add_4;             // value of pc + 4
    wire    [31: 0] NPC;            // next status of pc 
    wire    [31: 0] ExtOut;         // extention of 16-bit   
    wire    [31: 0] Ins;    // Ins gotten by im
    wire            Zero;           // zero generated by ALU

    wire    [31: 0] RegfileOut1;    // out1 of regfile
    wire    [31: 0] RegfileOut2;    // out2 of regfile

    wire    [ 4: 0] mux_RegDst_out;     // IM RF
    wire    [31: 0] mux_ALUSrc_out;    // RF ALU
    wire    [31: 0] mux_MemToReg_out;       // DM OUT

    wire    [3: 0] AluCtrlOut;     // out of alu controller
    wire    [31: 0] AluOut;         // out of alu
    wire    [31: 0] DmOut;          // out of dm
    wire    [31: 0] BeqPCOut;       // out of beq pc add 
    
    // DATAPATH
    pc pc(
        .clk(clk),
        .rst(rst),
        .PC(PC),
        .NPC(NPC)
    );

    PC_add pc_add4(
        .PC(PC),
        .PC_add_4(PC_add_4)
    );

    npc npc(
        .PC_add_4(PC_add_4), 
        .Branch(MEM_Branch),
        .Zero(MEM_Zero),
        .Jump(MEM_Jump),
        .Beq_ext_imm(MEM_Extimm),
        .Jump_ins_add(MEM_Jump_ins_add),
        .NPC(NPC)
    );

    im im(
        .PC(PC),
        .out_ins(Ins)
    );

    IF_ID IF_ID(
        .clk(clk),
        .IF_PC(PC_add_4),
        .IF_ins(Ins),

        .ID_PC(ID_PC),
        .ID_ins(ID_ins)
    );

    register_file register_files(
        .rs(ID_ins[25:21]),
        .rt(ID_ins[20:16]),
        .rd(WB_Reg_Write),
        .writedata(mux_MemToReg_out),
        .RegWrite(WB_RegWrite),
        .clk(clk),
        .rst(rst),

        .ReadData1(RegfileOut1),
        .ReadData2(RegfileOut2)
    );

    ID_EX ID_EX(
        .clk(clk),
        .ID_MemtoReg(MemtoReg),
        .ID_RegWrite(RegWrite),
        .ID_Branch(Branch),
        .ID_Jump(Jump),
        .ID_MemWrite(MemWrite),
        .ID_MemRead(MemRead),
        .ID_RegDst(RegDst),
        .ID_ALUSrc(ALUSrc),
        .ID_ExtOp(ExtOp),
        .ID_ALUOp(ALUOp),
        .ID_PC(ID_PC),
        .ID_Jump_ins_add(ID_ins[25:0]),
        .ID_ReadData1(RegfileOut1),
        .ID_ReadData2(RegfileOut2),
        .ID_Extimm(ID_ins[15:0]),
        .ID_rt(ID_ins[20:16]),
        .ID_rd(ID_ins[15:11]),

        .EX_MemtoReg(EX_MemtoReg),
        .EX_RegWrite(EX_RegWrite),
        .EX_Branch(EX_Branch),
        .EX_Jump(EX_Jump),
        .EX_MemWrite(EX_MemWrite),
        .EX_MemRead(EX_MemRead),
        .EX_RegDst(EX_RegDst),
        .EX_ALUSrc(EX_ALUSrc),
        .EX_ExtOp(EX_ExtOp),
        .EX_ALUOp(EX_ALUOp),
        .EX_PC(EX_PC),
        .EX_Jump_ins_add(EX_Jump_ins_add),
        .EX_ReadData1(EX_Reg_data_1_out),
        .EX_ReadData2(EX_Reg_data_2_out),
        .EX_Extimm(EX_Extimm),
        .EX_rt(EX_rt),
        .EX_rd(EX_rd)
    );

    mux_RegDst IF_ID_MUX(
        .rt(EX_rt),
        .rd(EX_rd),
        .RegDst(EX_RegDst),
        .mux_RegDst_out(mux_RegDst_out)
    );

    ext extend_immediate(
        .ins16(EX_Extimm),
        .ExtOp(EX_ExtOp),
        .Extimm(ExtOut)
    );

    mux_ALUSrc RF_ALU_MUX(
        .rtData(EX_Reg_data_2_out),
        .Imm(ExtOut),
        .ALUSrc(EX_ALUSrc),
        .mux_ALUSrc_out(mux_ALUSrc_out)
    );

    alu_ctrl ALU_controller(
        .func(ExtOut[5:0]),
        .ALUOp(EX_ALUOp),
        .AluCtrlOut(AluCtrlOut)
    );

    alu ALU(
        .rs(EX_Reg_data_1_out),
        .rt(mux_ALUSrc_out),
        .AluCtrlOut(AluCtrlOut),
        .Zero(Zero),
        .AluOut(AluOut)
    );

    EX_MEM EX_MEM(
        .clk(clk),
        .EX_MemtoReg(EX_MemtoReg),
        .EX_RegWrite(EX_RegWrite),
        .EX_Branch(EX_Branch),
        .EX_Jump(EX_Jump),
        .EX_MemWrite(EX_MemWrite),
        .EX_MemRead(EX_MemRead),
        .EX_PC(EX_PC),
        .EX_Jump_ins_add(EX_Jump_ins_add),
        .EX_Zero(Zero),
        .EX_ALU(AluOut),
        .EX_WriteData(EX_Reg_data_2_out),
        .EX_Extimm(ExtOut),
        .EX_Reg_Write(mux_RegDst_out),

        .MEM_MemtoReg(MEM_MemtoReg),
        .MEM_RegWrite(MEM_RegWrite),
        .MEM_Branch(MEM_Branch),
        .MEM_Jump(MEM_Jump),
        .MEM_MemWrite(MEM_MemWrite),
        .MEM_MemRead(MEM_MemRead),
        .MEM_PC(MEM_PC),
        .MEM_Jump_ins_add(MEM_Jump_ins_add),
        .MEM_Zero(MEM_Zero),
        .MEM_ALU(MEM_ALU),
        .MEM_WriteData(MEM_WriteData),
        .MEM_Extimm(MEM_Extimm),
        .MEM_Reg_Write(MEM_Reg_Write)
    );

    dm data_memory(
        .MEM_ALU(MEM_ALU),
        .MEM_WriteData(MEM_WriteData),
        .MemWrite(MEM_MemWrite),
        .MemRead(MEM_MemRead),
        .clk(clk),

        .dm_out(DmOut)
    );

    MEM_WB MEM_WB(
        .clk(clk),
        .MEM_MemtoReg(MEM_MemtoReg),
        .MEM_RegWrite(MEM_RegWrite),
        .MEM_Data_in(DmOut),
        .MEM_ALU(MEM_ALU),
        .MEM_Reg_Write(MEM_Reg_Write),

        .WB_MemtoReg(WB_MemtoReg),
        .WB_RegWrite(WB_RegWrite),
        .WB_Data_out(WB_Data_out),
        .WB_ALU(WB_ALU),
        .WB_Reg_Write(WB_Reg_Write)
    );

    mux_MemToReg DM_OUT_MUX(
        .DmData(WB_Data_out),
        .ALUData(WB_ALU),
        .MemtoReg(WB_MemtoReg),

        .mux_MemToReg_out(mux_MemToReg_out)
    );
endmodule //data_path
