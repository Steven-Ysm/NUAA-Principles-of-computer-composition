`include "./controller/ctrl.v"

`include "./datapath/alu_ctrl.v"
`include "./datapath/alu.v"
`include "./datapath/dm.v"
`include "./datapath/Ext.v"
`include "./datapath/im.v"
`include "./datapath/mux.v"
`include "./datapath/npc.v"
`include "./datapath/pc.v"
`include "./datapath/registerfile.v"

`include "./datapath/EX_MEM.v"
`include "./datapath/ID_EX.v"
`include "./datapath/IF_ID.v"
`include "./datapath/MEM_WB.v"

`include "./datapath/hazard_and_forward.v"
`include "./datapath/compare.v"

module Mips(clk,rst);

    input clk;
    input rst;

    wire RegDst;
    wire Branch;
    wire MemtoReg;
    wire MemWrite;
    wire ALUSrc;
    wire RegWrite;
    wire Jump;
    wire Ext_op;

    wire [2:0] ALUOp;

    wire [31:0] instruction;

    wire [31:0] PC; 
    wire [31:0] NPC; 
    wire [31:0] ext_out;   
    wire zero; // zero generated by ALU

    wire [31:0] regfile_out1; 
    wire [31:0] regfile_out2; 

    wire [4:0] mux_RegDst_out;
    wire [31:0] mux_ALUSrc_out; 
    wire [31:0] mux_MemToReg_out;

    wire [2:0] alu_ctrl_out; 
    wire [31:0] alu_out; 
    wire [31:0] dm_out; 
    wire undefine;
    wire overflow;

    //if_id
    wire [31:0] ID_ins;
    wire [31:0] ID_PC;

    //id_ex
    wire EX_RegDst;   
    wire EX_Branch;
    wire EX_MemtoReg;
    wire EX_MemWrite;
    wire EX_ALUSrc;
    wire EX_RegWrite;
    wire EX_Jump;
    wire EX_Ext_op;  
    wire [31:0]  EX_ReadData1;
    wire [31:0]  EX_ReadData2;
    wire [31:0]  EX_PC;
    wire [25:0]  EX_ins;
    wire [2:0] EX_ALUOp;

    //ex_mem          
    wire MEM_Branch;
    wire MEM_Jump;
    wire MEM_MemtoReg;
    wire MEM_MemWrite;
    wire MEM_RegWrite;
    wire MEM_zero;
    wire MEM_undefine;

    wire [25:0] MEM_jump_Addr;
    wire [31:0] PC_Branch;
    wire [31:0] MEM_pc;
    wire [31:0] MEM_alu_out;
    wire [31:0] MEM_ReadData2;
    wire [4:0] MEM_mux_RegDst_out;

    //mem_wb
    wire WB_MemtoReg;
    wire WB_RegWrite;
    
    wire [31:0] WB_dm_out;
    wire [31:0] WB_alu_out;
    wire [4:0] rd;

    //hazard && forward
    wire PCWrite;
    wire IFWrite;
    wire flushE;
    wire IFflush;

    wire [31:0] mux_forward_out_1;
    wire [31:0] mux_forward_out_2;
    
    //Forward
    wire Compare_Zero;
    wire [1:0] forwardrs;
    wire [1:0] forwardrt;
    wire [1:0] forwardrsd;             
    wire [1:0] forwardrtd;
    
    wire [31:0] EX_Extimm;

    pc pc(
        .clk(clk),
        .rst(rst),
        .NPC(NPC),
        .PC(PC),
        .PCWrite(PCWrite)
    );

    npc npc(
        .PC(PC),
        .Branch(Branch),
        .Compare_Zero(Compare_Zero),
        .Jump(Jump),
        .PC_add_4(ID_PC),
        .Beq_ext_imm(ext_out),
        .Jump_ins_add(ID_ins),
        .NPC(NPC)
    );

    im im(
        .PC(PC),
        .out_ins(instruction)
    );

    IF_ID if_id(
        .clk(clk),
        .rst(rst),

        .IF_ins(instruction),
        .ID_ins(ID_ins),
        .IF_PC(PC),
        .ID_PC(ID_PC),
        
        .IFWrite(IFWrite),
        .IFflush(IFflush)
    );

    ctrl Ctrl(
        .Opcode(ID_ins[31:26]),
        .RegDst(RegDst),
        .Branch(Branch),
        .MemtoReg(MemtoReg),
        .ALUOp(ALUOp),
        .MemWrite(MemWrite),
        .ALUSrc(ALUSrc),
        .RegWrite(RegWrite),
        .Jump(Jump),
        .Ext_op(Ext_op)
    );

    mux_RegDst IF_ID_MUX(
        .rt(EX_ins[20:16]),
        .rd(EX_ins[15:11]),
        .EX_RegDst(EX_RegDst),
        .mux_RegDst_out(mux_RegDst_out)
    );

    register_file register_files(
        .rs(ID_ins[25:21]),
        .rt(ID_ins[20:16]),
        .rd(rd),
        .writedata(mux_MemToReg_out),
        .WB_RegWrite(WB_RegWrite),
        .clk(clk),
        .rst(rst),
        .ReadData1(regfile_out1),
        .ReadData2(regfile_out2)
    );

    ID_EX idex(
        .clk(clk),
        .rst(rst),
        .EXflush(flushE),

        .ReadData1(regfile_out1),
        .ReadData2(regfile_out2),
        .ID_PC(ID_PC),
        .ID_ins(ID_ins[25:0]),
        .Extimm(ext_out),
        
        .RegDst(RegDst),
        .Branch(Branch),
        .MemtoReg(MemtoReg), 
        .ALUOp(ALUOp), 
        .MemWrite(MemWrite), 
        .ALUSrc(ALUSrc), 
        .RegWrite(RegWrite), 
        .Jump(Jump), 
        .Ext_op(Ext_op),
        

        .EX_ReadData1(EX_ReadData1),
        .EX_ReadData2(EX_ReadData2),
        .EX_ins(EX_ins),
        .EX_PC(EX_PC),
        .EX_Extimm(EX_Extimm),

        .EX_RegDst(EX_RegDst),
        .EX_Branch(EX_Branch),
        .EX_MemtoReg(EX_MemtoReg),
        .EX_ALUOp(EX_ALUOp),
        .EX_MemWrite(EX_MemWrite),
        .EX_ALUSrc(EX_ALUSrc),
        .EX_RegWrite(EX_RegWrite),
        .EX_Jump(EX_Jump),
        .EX_Ext_op(EX_Ext_op)
    );

    mux_forward Forward_MUX_1(
        .forward(forwardrs),
        .EX_ReadData(EX_ReadData1),
        .mux_MemToReg_out(mux_MemToReg_out),
        .MEM_AluOut(MEM_alu_out),

        .mux_forward_out(mux_forward_out_1)
    );


    mux_forward Forward_MUX_2(
        .forward(forwardrt),
        .EX_ReadData(EX_ReadData2),
        .mux_MemToReg_out(mux_MemToReg_out),
        .MEM_AluOut(MEM_alu_out),

        .mux_forward_out(mux_forward_out_2)
    );

    Ext extension_unit(
        .ins16(ID_ins[15:0]),
        .Ext_op(Ext_op),
        .Extimm(ext_out) 
    );

    mux_ALUSrc RF_ALU_MUX(
        .mux_forward_out2(mux_forward_out_2),
        .Extimm(EX_Extimm),
        .EX_ALUSrc(EX_ALUSrc),
        .mux_ALUSrc_out(mux_ALUSrc_out)
    );

    alu_ctrl ALU_controller(
        .func(EX_ins[5:0]),
        .EX_ALUOp(EX_ALUOp),
        .AluCtrlOut(alu_ctrl_out),
        .undefine(undefine)
    );

    alu ALU(
        .A(mux_forward_out_1),
        .B(mux_ALUSrc_out),
        .AluCtrlOut(alu_ctrl_out),
        .zero(zero),
        .AluOut(alu_out),
        .overflow(overflow)
    );

    EX_MEM exmem(
        .clk(clk),
        .rst(rst),

        .EX_PC(EX_PC),
        .EX_ins(EX_ins),
        .Extimm(ext_out),
        .AluOut(alu_out),
        .EX_ReadData2(EX_ReadData2),
        .mux_RegDst_out(mux_RegDst_out),

        .EX_Branch(EX_Branch), 
        .EX_MemtoReg(EX_MemtoReg), 
        .EX_MemWrite(EX_MemWrite), 
        .EX_RegWrite(EX_RegWrite), 
        .EX_Jump(EX_Jump),

        .zero(zero),
        .undefine(undefine),
        .overflow(overflow),

        .MEM_PC(MEM_pc),
        .Jump_Addr(MEM_jump_Addr),
        .PC_Branch(PC_Branch),
        .MEM_AluOut(MEM_alu_out),
        .MEM_ReadData2(MEM_ReadData2),
        .MEM_mux_RegDst_out(MEM_mux_RegDst_out),

        .MEM_Branch(MEM_Branch),
        .MEM_MemtoReg(MEM_MemtoReg),
        .MEM_MemWrite(MEM_MemWrite),
        .MEM_RegWrite(MEM_RegWrite),
        .MEM_Jump(MEM_Jump),
    
        .MEM_zero(MEM_zero),
        .MEM_undefine(MEM_undefine),
        .MEM_overflow(MEM_overflow)
    );

    dm_4k data_memory(
        .clk(clk),
        .MEM_MemWrite(MEM_MemWrite),

        .MEM_AluOut(MEM_alu_out),
        .MEM_writedata(MEM_ReadData2),
        
        .dm_out(dm_out)
    );

    MEM_WB memwb(
        .clk(clk),
        .rst(rst),
        .MEM_MemtoReg(MEM_MemtoReg),
        .MEM_RegWrite(MEM_RegWrite),

        .dm_out(dm_out),
        .MEM_AluOut(MEM_alu_out),
        .MEM_mux_RegDst_out(MEM_mux_RegDst_out),
        .MEM_PC(MEM_pc),
        .MEM_undefine(MEM_undefine),
        .MEM_overflow(MEM_overflow),

        .WB_MemtoReg(WB_MemtoReg),
        .WB_RegWrite(WB_RegWrite),
        .WB_dm_out(WB_dm_out),
        .WB_AluOut(WB_alu_out),
        .rd(rd)
    );



    mux_MemToReg DM_OUT_MUX(
        .WB_dm_out(WB_dm_out),
        .WB_AluOut(WB_alu_out),
        .WB_MemtoReg(WB_MemtoReg),
        .mux_MemToReg_out(mux_MemToReg_out)
    );

    Hazard_and_Forward hazd_forward(
        .MEM_RegWrite(MEM_RegWrite),
        .MEM_MemtoReg(MEM_MemtoReg),
        .WB_RegWrite(WB_RegWrite),
        .Compare_Zero(Compare_Zero),

        .MEM_mux_RegDst_out(MEM_mux_RegDst_out),
        .rd(rd),
        .EX_rs(EX_ins[25:21]),
        .EX_rt(EX_ins[20:16]),
        .ID_rs(ID_ins[25:21]),
        .ID_rt(ID_ins[20:16]),
        .mux_RegDst_out(mux_RegDst_out),

        .forwardrs(forwardrs),
        .forwardrt(forwardrt),
        .PCWrite(PCWrite),
        .IFWrite(IFWrite),
        .EXflush(flushE),

        .Jump(Jump),
        .Branch(Branch),
        .EX_RegWrite(EX_RegWrite),
        .EX_MemtoReg(EX_MemtoReg),
        .EX_MemWrite(EX_MemWrite),
        
        .forward_rs_compare(forwardrsd),
        .forward_rt_compare(forwardrtd),
        .IFflush(IFflush)
    );
    
    Compare compare(
        .ReadData1(regfile_out1),
        .MEM_AluOut(MEM_alu_out),
        .forwardrsd(forwardrsd),
        
        .ReadData2(regfile_out2),
        .forwardrtd(forwardrtd),
        .AluOut(alu_out),

        .Compare_Zero(Compare_Zero)
    );

endmodule